// Code your design here
`include "dassign3.v"