// Code your testbench here
// or browse Examples
`include "dassign3.tb.v"